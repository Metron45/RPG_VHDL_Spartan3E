----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:22:56 05/07/2019 
-- Design Name: 
-- Module Name:    GameLogic - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity GameLogic is
   Port(
           DIV_X : in  STD_LOGIC_VECTOR (4 downto 0);
           DIV_Y : in  STD_LOGIC_VECTOR (3 downto 0);
           RGB_MAP : out  STD_LOGIC_VECTOR (2 downto 0) 
       );
end GameLogic;

architecture Behavioral of GameLogic is
signal x: integer range 0 to 20;
signal y: integer range 0 to 15;
type ARRAY_2D is array ( (20*15) -1 downto 0) of std_logic_vector (2 downto 0);
constant Territory : ARRAY_2D := (  "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101",
                                    "000", "001", "010", "011", "100", "101", "110", "111", "101", "010",
                                    "010", "000", "001", "010", "011", "100", "101", "110", "111", "101"  );

begin
x <= to_integer( unsigned( DIV_X ) );
y <= to_integer( unsigned( DIV_Y ) );

process(x,y)
begin
   RGB_MAP <= Territory( y*4 + x );
end process;

end Behavioral;

